module top
    (
        
    );


endmodule
