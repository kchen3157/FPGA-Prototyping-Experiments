

module sseg
endmodule